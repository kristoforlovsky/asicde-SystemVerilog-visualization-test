module TestModule (
);


Mod1 1 (
  .I1    (),
  .I2    (),
  .O1    (),
  .O2    ()
);


endmodule: TestModule